LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.all;

entity datapath is
	port(clk: in std_logic
	);
end datapath;

architecture arch of datapath is
	
		
		
end arch;